// crypto IP

module crypto (
  input logic [99:0] a,
  input logic [99:0] b,
  input logic clk,
  output logic [99:0] out
);

  wire [99:0] clk_skew;
  
endmodule
